library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.ALL;

entity instr_mem is
	generic(
		operand_width : integer:=16
        );
	port (
		mem_add: in std_logic_vector((operand_width - 1) downto 0);
        mem_data: out std_logic_vector((operand_width - 1) downto 0)
        );
end instr_mem;

architecture behavioural of instr_mem is
    type memm is array (0 to 127) of std_logic_vector((operand_width - 1) downto 0);
	 signal sData: memm := (others => (others => '0'));
begin
    mem_read: process(mem_add)
        variable Data: memm := (
	     0 => "0001001010011000", -- ADD
	     1 => "0001001010011011", 
	     2 => "0001001010011000", 
	     3 => "0001001010011011", 
	     4 => "0001001010011000", 
	     5 => "0001001010011011", 
	     6 => "0001001010011000", 
	     7 => "0011001000000000", --LLI R1 0
	     8 => "0011010000000000", --LLI R2 0
	     9 => "0011100000000111", --LLI R4 3
		 10 => "0001011110111000", --ADA R3,R6,R7
	    11 => "0011001000000001", 
	    12 => "0011010000000010", 
	    13 => "0011001000000011", 
	    14 => "0011010000000100", 
	    15 => "0011001000000101", 		 
	    16 => "0011010000000000", 		 
		 --17 => "0001111011100001",	--ADZ R7,R3,R4		
		 --17 => "0100110100000000",	--LW R6, R4,0 	    
		 --17 => "0101100011000010", --SW R4,R3,2
		 17 =>
		 18 => "0011001000000001", 
	    19 => "0011010000000010", 
	    20 => "0011001000000011", 
	    21 => "0011010000000100", 
	    22 => "0011001000000101", 		 
	    23 => "0011010000000110", 		  
	    24 => "0011010000000111", 
	    25 => "0011001000001000", 	 
		 26 => "0100110111000010s",	--LW R6, R4,0 	
	    27 => "0011001000000011", 
	    28 => "0011010000000100", 
	    29 => "0011001000000101",  
	    30 => "0011010000000110",   
	    31 => "0011010000000111", 
	    32 => "0011001000001000", 
		 33 => "0000111100000110", 	 
	    34 => "0011001000000011", 
	    35 => "0011010000000100", 
	    36 => "0011001000000101", 		 
	    37 => "0011010000000110", 		  
	    38 => "0011010000000111", 
	    39 => "0011001000001000", 		 

		 
	     others => (others => '0')
	 );
	 begin
    mem_data <= Data(to_integer(unsigned(mem_add)));
	 sData <= Data;
    end process;
end architecture;